module top_cpu #(
    parameter WORD_WIDTH = 32,     //字长
    parameter ADDR_WIDTH = 32      //地址宽度
)(
    input clk,
    input rstn,
    input rxd,
    output txd
);
    












endmodule