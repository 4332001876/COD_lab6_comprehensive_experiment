module cache_direct_mapped(

);







endmodule